localparam [5:0]IP_pos[0:63] = {
	57,49,41,33,25,17,9,1, 
	59,51,43,35,27,19,11,3, 
	61,53,45,37,29,21,13,5, 
	63,55,47,39,31,23,15,7, 
	56,48,40,32,24,16,8,0, 
	58,50,42,34,26,18,10,2, 
	60,52,44,36,28,20,12,4, 
	62,54,46,38,30,22,14,6
};

localparam [4:0]E_pos[0:47] = {
	31,0,1,2,3,4,
	3,4,5,6,7,8,
	7,8,9,10,11,12,
	11,12,13,14,15,16,
	15,16,17,18,19,20,
	19,20,21,22,23,24,
	23,24,25,26,27,28,
	27,28,29,30,31,0
};

localparam [4:0]P_pos[0:31] = {
	15,6,19,20, 
	28,11,27,16, 
	0,14,22,25, 
	4,17,30,9, 
	1,7,23,13, 
	31,26,2,8, 
	18,12,29,5, 
	21,10,3,24
};

localparam [6:0]PC1_pos[0:55] = {
	56,48,40,32,24,16,8, 
	0,57,49,41,33,25,17, 
	9,1,58,50,42,34,26, 
	18,10,2,59,51,43,35, 
	62,54,46,38,30,22,14, 
	6,61,53,45,37,29,21, 
	13,5,60,52,44,36,28, 
	20,12,4,27,19,11,3
};

localparam [5:0]PC2_pos[0:47] = {
	13,16,10,23,0,4,
	2,27,14,5,20,9,
	22,18,11,3,25,7,
	15,6,26,19,12,1,
	40,51,30,36,46,54,
	29,39,50,44,32,47,
	43,48,38,55,33,52,
	45,41,49,35,28,31
};

localparam [5:0]IP_inv_pos[0:63] = {
	39,7,47,15,55,23,63,31, 
	38,6,46,14,54,22,62,30, 
	37,5,45,13,53,21,61,29, 
	36,4,44,12,52,20,60,28, 
	35,3,43,11,51,19,59,27, 
	34,2,42,10,50,18,58,26, 
	33,1,41,9,49,17,57,25, 
	32,0,40,8,48,16,56,24
};

localparam [3:0]S_val[0:7][0:63] = '{ '{
	14, 4, 13, 1, 2, 15, 11, 8, 3, 10, 6, 12, 5, 9, 0, 7, 
	0, 15, 7, 4, 14, 2, 13, 1, 10, 6, 12, 11, 9, 5, 3, 8, 
	4, 1, 14, 8, 13, 6, 2, 11, 15, 12, 9, 7, 3, 10, 5, 0, 
	15, 12, 8, 2, 4, 9, 1, 7, 5, 11, 3, 14, 10, 0, 6, 13
},'{
	15, 1, 8, 14, 6, 11, 3, 4, 9, 7, 2, 13, 12, 0, 5, 10, 
	3, 13, 4, 7, 15, 2, 8, 14, 12, 0, 1, 10, 6, 9, 11, 5, 
	0, 14, 7, 11, 10, 4, 13, 1, 5, 8, 12, 6, 9, 3, 2, 15, 
	13, 8, 10, 1, 3, 15, 4, 2, 11, 6, 7, 12, 0, 5, 14, 9
},'{
	10, 0, 9, 14, 6, 3, 15, 5, 1, 13, 12, 7, 11, 4, 2, 8, 
	13, 7, 0, 9, 3, 4, 6, 10, 2, 8, 5, 14, 12, 11, 15, 1, 
	13, 6, 4, 9, 8, 15, 3, 0, 11, 1, 2, 12, 5, 10, 14, 7, 
	1, 10, 13, 0, 6, 9, 8, 7, 4, 15, 14, 3, 11, 5, 2, 12
},'{
	7, 13, 14, 3, 0, 6, 9, 10, 1, 2, 8, 5, 11, 12, 4, 15, 
	13, 8, 11, 5, 6, 15, 0, 3, 4, 7, 2, 12, 1, 10, 14, 9, 
	10, 6, 9, 0, 12, 11, 7, 13, 15, 1, 3, 14, 5, 2, 8, 4, 
	3, 15, 0, 6, 10, 1, 13, 8, 9, 4, 5, 11, 12, 7, 2, 14
},'{
	2, 12, 4, 1, 7, 10, 11, 6, 8, 5, 3, 15, 13, 0, 14, 9, 
	14, 11, 2, 12, 4, 7, 13, 1, 5, 0, 15, 10, 3, 9, 8, 6, 
	4, 2, 1, 11, 10, 13, 7, 8, 15, 9, 12, 5, 6, 3, 0, 14, 
	11, 8, 12, 7, 1, 14, 2, 13, 6, 15, 0, 9, 10, 4, 5, 3
},'{
	12, 1, 10, 15, 9, 2, 6, 8, 0, 13, 3, 4, 14, 7, 5, 11, 
	10, 15, 4, 2, 7, 12, 9, 5, 6, 1, 13, 14, 0, 11, 3, 8, 
	9, 14, 15, 5, 2, 8, 12, 3, 7, 0, 4, 10, 1, 13, 11, 6, 
	4, 3, 2, 12, 9, 5, 15, 10, 11, 14, 1, 7, 6, 0, 8, 13
},'{
	4, 11, 2, 14, 15, 0, 8, 13, 3, 12, 9, 7, 5, 10, 6, 1, 
	13, 0, 11, 7, 4, 9, 1, 10, 14, 3, 5, 12, 2, 15, 8, 6, 
	1, 4, 11, 13, 12, 3, 7, 14, 10, 15, 6, 8, 0, 5, 9, 2, 
	6, 11, 13, 8, 1, 4, 10, 7, 9, 5, 0, 15, 14, 2, 3, 12
},'{
	13, 2, 8, 4, 6, 15, 11, 1, 10, 9, 3, 14, 5, 0, 12, 7, 
	1, 15, 13, 8, 10, 3, 7, 4, 12, 5, 6, 11, 0, 14, 9, 2, 
	7, 11, 4, 1, 9, 12, 14, 2, 0, 6, 10, 13, 15, 3, 5, 8, 
	2, 1, 14, 7, 4, 10, 8, 13, 15, 12, 9, 0, 3, 5, 6, 11
} };


function [0:63]IP(input [0:63] in);
	for(int i = 0; i < 64; i++) IP[i] = in[IP_pos[i]];
endfunction

function [0:47]E(input [0:31] in);
	for(int i = 0; i < 48; i++) E[i] = in[E_pos[i]];
endfunction

function [0:31]P(input [0:31] in);
	for(int i = 0; i < 32; i++) P[i] = in[P_pos[i]];
endfunction

function [0:55]PC1(input [0:63] in);
	for(int i = 0; i < 56; i++) PC1[i] = in[PC1_pos[i]];
endfunction

function [0:47]PC2(input [0:55] in);
	for(int i = 0; i < 48; i++) PC2[i] = in[PC2_pos[i]];
endfunction

function [0:63]IP_inv(input [0:63] in);
	for(int i = 0; i < 64; i++) IP_inv[i] = in[IP_inv_pos[i]];
endfunction

function [0:31]S(input[0:47] in);
	for(int i = 0; i < 8; i++) S[i*4 +: 4] = S_val[i][ ({in[i*6], in[(i*6)+5]} * 16) + in[(i*6)+1 +: 4] ];
endfunction

function [0:63]DES_round(input[0:63] in, input[0:47] k);
	DES_round[0:31] = in[32:63];
	DES_round[32:63] = in[0:31] ^ P( S( E( in[32:63] ) ^ k ) );
endfunction

function count_to_shift_n(input [3:0] cnt);
	casez(cnt)
		4'd0, 4'd1, 4'd8, 4'd15 : count_to_shift_n = 1'b0;
		default                   count_to_shift_n = 1'b1;
	endcase
endfunction

function automatic[0:55]DES_key_cd_shift(
	input[0:55] in, 
	input dir, 		// deasserted shift left, asserted shift right
	input n			// deasserted shift 1, asserted shift 2
);
	logic  [0:27] c = in[0:27];
	logic  [0:27] d = in[28:55];

	casez({dir,n})
		2'b00 : DES_key_cd_shift = {c[1:27], c[0],      d[1:27], d[0]};
		2'b01 : DES_key_cd_shift = {c[2:27], c[0:1],    d[2:27], d[0:1]};
		2'b10 : DES_key_cd_shift = {c[27], c[0:26],     d[27], d[0:26]};
		2'b11 : DES_key_cd_shift = {c[26:27], c[0:25],  d[26:27], d[0:25]};
	endcase
endfunction
